`timescale 1ns / 1ps

module font_rom(
    input  wire        clk,
    input  wire [7:0]  char_code,   // ex: '0', '1', '+', '=' ASCII
    input  wire [3:0]  row,         // 0~7 row (y-direction)
    output reg  [7:0]  font_line    // 8 pixels in one row (x-direction)
);

    reg [7:0] rom [0:127][0:7]; // 128 ASCII chars, 8 rows each

    initial begin
        // Digits '0' to '9'
        rom[8'd48][0] = 8'b00111100;
        rom[8'd48][1] = 8'b01100110;
        rom[8'd48][2] = 8'b01101110;
        rom[8'd48][3] = 8'b01110110;
        rom[8'd48][4] = 8'b01100110;
        rom[8'd48][5] = 8'b01100110;
        rom[8'd48][6] = 8'b00111100;
        rom[8'd48][7] = 8'b00000000;

        rom[8'd49][0] = 8'b00011000;
        rom[8'd49][1] = 8'b00111000;
        rom[8'd49][2] = 8'b00011000;
        rom[8'd49][3] = 8'b00011000;
        rom[8'd49][4] = 8'b00011000;
        rom[8'd49][5] = 8'b00011000;
        rom[8'd49][6] = 8'b00111100;
        rom[8'd49][7] = 8'b00000000;

        rom[8'd50][0] = 8'b00111100;
        rom[8'd50][1] = 8'b01100110;
        rom[8'd50][2] = 8'b00000110;
        rom[8'd50][3] = 8'b00001100;
        rom[8'd50][4] = 8'b00110000;
        rom[8'd50][5] = 8'b01100000;
        rom[8'd50][6] = 8'b01111110;
        rom[8'd50][7] = 8'b00000000;

        rom[8'd51][0] = 8'b00111100;
        rom[8'd51][1] = 8'b01100110;
        rom[8'd51][2] = 8'b00000110;
        rom[8'd51][3] = 8'b00011100;
        rom[8'd51][4] = 8'b00000110;
        rom[8'd51][5] = 8'b01100110;
        rom[8'd51][6] = 8'b00111100;
        rom[8'd51][7] = 8'b00000000;

        rom[8'd52][0] = 8'b00001100;
        rom[8'd52][1] = 8'b00011100;
        rom[8'd52][2] = 8'b00111100;
        rom[8'd52][3] = 8'b01101100;
        rom[8'd52][4] = 8'b01111110;
        rom[8'd52][5] = 8'b00001100;
        rom[8'd52][6] = 8'b00011110;
        rom[8'd52][7] = 8'b00000000;

        rom[8'd53][0] = 8'b01111110;
        rom[8'd53][1] = 8'b01100000;
        rom[8'd53][2] = 8'b01111100;
        rom[8'd53][3] = 8'b00000110;
        rom[8'd53][4] = 8'b00000110;
        rom[8'd53][5] = 8'b01100110;
        rom[8'd53][6] = 8'b00111100;
        rom[8'd53][7] = 8'b00000000;

        rom[8'd54][0] = 8'b00111100;
        rom[8'd54][1] = 8'b01100110;
        rom[8'd54][2] = 8'b01100000;
        rom[8'd54][3] = 8'b01111100;
        rom[8'd54][4] = 8'b01100110;
        rom[8'd54][5] = 8'b01100110;
        rom[8'd54][6] = 8'b00111100;
        rom[8'd54][7] = 8'b00000000;

        rom[8'd55][0] = 8'b01111110;
        rom[8'd55][1] = 8'b00000110;
        rom[8'd55][2] = 8'b00001100;
        rom[8'd55][3] = 8'b00011000;
        rom[8'd55][4] = 8'b00110000;
        rom[8'd55][5] = 8'b00110000;
        rom[8'd55][6] = 8'b00110000;
        rom[8'd55][7] = 8'b00000000;

        rom[8'd56][0] = 8'b00111100;
        rom[8'd56][1] = 8'b01100110;
        rom[8'd56][2] = 8'b01100110;
        rom[8'd56][3] = 8'b00111100;
        rom[8'd56][4] = 8'b01100110;
        rom[8'd56][5] = 8'b01100110;
        rom[8'd56][6] = 8'b00111100;
        rom[8'd56][7] = 8'b00000000;

        rom[8'd57][0] = 8'b00111100;
        rom[8'd57][1] = 8'b01100110;
        rom[8'd57][2] = 8'b01100110;
        rom[8'd57][3] = 8'b00111110;
        rom[8'd57][4] = 8'b00000110;
        rom[8'd57][5] = 8'b01100110;
        rom[8'd57][6] = 8'b00111100;
        rom[8'd57][7] = 8'b00000000;

        // '+' symbol (ASCII 43)
        rom[8'd43][0] = 8'b00011000;
        rom[8'd43][1] = 8'b00011000;
        rom[8'd43][2] = 8'b00011000;
        rom[8'd43][3] = 8'b11111111;
        rom[8'd43][4] = 8'b00011000;
        rom[8'd43][5] = 8'b00011000;
        rom[8'd43][6] = 8'b00011000;
        rom[8'd43][7] = 8'b00000000;

        // '=' symbol (ASCII 61)
        rom[8'd61][0] = 8'b00000000;
        rom[8'd61][1] = 8'b11111111;
        rom[8'd61][2] = 8'b00000000;
        rom[8'd61][3] = 8'b00000000;
        rom[8'd61][4] = 8'b11111111;
        rom[8'd61][5] = 8'b00000000;
        rom[8'd61][6] = 8'b00000000;
        rom[8'd61][7] = 8'b00000000;
    end

    always @(posedge clk)
        font_line <= rom[char_code][row];

endmodule
